interface rx_intf;
logic rx_tlast_i;
logic rx_tvalid_i;
logic [15:0]rx_tdata_i;

logic rx_tready_o;

logic aclk_i;
logic aresetn_i;


endinterface
