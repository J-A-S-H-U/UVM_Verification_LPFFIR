package top_pkg;

	import uvm_pkg::*
	`include "uvm_macros.svh"
	
	import rx_pkg.sv::*;
	import tx_pkg.sv::*;
	
	`include "reference.sv"
	`include "scoreboard.sv"
	`include "environment.sv"
	`include "test.sv"
endpackage