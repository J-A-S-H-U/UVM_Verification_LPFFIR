package rx_pkg;

	import uvm_pkg::*
	`include "uvm_macros.svh"
	
	`include "rx_intf.sv"
	`include "rx_seq_item.sv"
	`include "rx_sequence.sv"
	`include "rx_sequencer.sv"
	`include "rx_driver.sv"
	`include "rx_monitor.sv"
	`include "rx_agent.sv"
endpackage