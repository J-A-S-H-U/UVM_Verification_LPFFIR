interface tx_intf;
logic tx_tlast_o;
logic tx_tvalid_o;
logic [15:0]tx_tdata_o;

logic tx_tready_i;

logic aclk_i;
logic aresetn_i;


endinterface