package tx_pkg;

	import uvm_pkg::*
	`include "uvm_macros.svh"
	
	`include "tx_intf.sv"
	`include "tx_seq_item.sv"
	`include "tx_sequence.sv"
	`include "tx_sequencer.sv"
	`include "tx_driver.sv"
	`include "tx_monitor.sv"
	`include "tx_agent.sv"
endpackage